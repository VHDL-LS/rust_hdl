-- Package env as defined by IEEE 1076-2008

package env is
end package;

-- Package texio as defined by IEEE 1076-2008

package textio is
end package;
